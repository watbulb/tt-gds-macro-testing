`ifndef BLACKBOX_NAME
`define BLACKBOX_NAME ttlogo
`endif
`ifndef BLACKBOX_INSTANCE
`define BLACKBOX_INSTANCE um_ttlogo
`endif

(* blackbox *) (* keep *)
module `BLACKBOX_NAME ();
endmodule

