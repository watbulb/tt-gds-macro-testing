`ifndef BLACKBOX_NAME
`define BLACKBOX_NAME skullfet_logo
`endif
`ifndef BLACKBOX_INSTANCE
`define BLACKBOX_INSTANCE um_skullfet_logo
`endif

(* blackbox *) (* keep *)
module `BLACKBOX_NAME ();
endmodule

