VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ttlogo
  CLASS BLOCK ;
  FOREIGN ttlogo ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 35.840 ;
  OBS
      LAYER met2 ;
        RECT 16.800 35.560 19.320 35.840 ;
        RECT 14.560 35.280 21.560 35.560 ;
        RECT 13.440 35.000 22.680 35.280 ;
        RECT 12.600 34.720 23.520 35.000 ;
        RECT 11.760 34.440 24.360 34.720 ;
        RECT 10.920 34.160 25.200 34.440 ;
        RECT 10.360 33.880 25.760 34.160 ;
        RECT 9.800 33.600 26.320 33.880 ;
        RECT 9.240 33.320 26.880 33.600 ;
        RECT 8.680 33.040 27.440 33.320 ;
        RECT 8.400 32.760 27.720 33.040 ;
        RECT 7.840 32.480 15.120 32.760 ;
        RECT 21.000 32.480 28.280 32.760 ;
        RECT 7.560 32.200 14.000 32.480 ;
        RECT 22.120 32.200 28.560 32.480 ;
        RECT 7.280 31.920 13.160 32.200 ;
        RECT 22.960 31.920 28.840 32.200 ;
        RECT 6.720 31.640 12.320 31.920 ;
        RECT 23.800 31.640 29.400 31.920 ;
        RECT 6.440 31.360 11.760 31.640 ;
        RECT 24.360 31.360 29.680 31.640 ;
        RECT 6.160 31.080 11.200 31.360 ;
        RECT 24.920 31.080 29.960 31.360 ;
        RECT 5.880 30.800 10.640 31.080 ;
        RECT 25.480 30.800 30.240 31.080 ;
        RECT 5.600 30.520 10.080 30.800 ;
        RECT 26.040 30.520 30.520 30.800 ;
        RECT 5.320 30.240 9.800 30.520 ;
        RECT 26.320 30.240 30.800 30.520 ;
        RECT 5.040 29.960 9.240 30.240 ;
        RECT 26.880 29.960 31.080 30.240 ;
        RECT 4.760 29.680 8.960 29.960 ;
        RECT 27.160 29.680 31.360 29.960 ;
        RECT 4.480 29.400 8.680 29.680 ;
        RECT 27.440 29.400 31.640 29.680 ;
        RECT 4.200 29.120 8.120 29.400 ;
        RECT 28.000 29.120 31.920 29.400 ;
        RECT 3.920 28.840 7.840 29.120 ;
        RECT 28.280 28.840 32.200 29.120 ;
        RECT 3.920 28.560 7.560 28.840 ;
        RECT 28.560 28.560 32.200 28.840 ;
        RECT 3.640 28.280 7.280 28.560 ;
        RECT 28.840 28.280 32.480 28.560 ;
        RECT 3.360 28.000 21.560 28.280 ;
        RECT 29.120 28.000 32.760 28.280 ;
        RECT 3.080 27.440 21.560 28.000 ;
        RECT 29.400 27.720 33.040 28.000 ;
        RECT 2.800 27.160 21.560 27.440 ;
        RECT 29.680 27.440 33.040 27.720 ;
        RECT 29.680 27.160 33.320 27.440 ;
        RECT 2.520 26.600 21.560 27.160 ;
        RECT 29.960 26.880 33.600 27.160 ;
        RECT 30.240 26.600 33.600 26.880 ;
        RECT 2.240 26.040 21.560 26.600 ;
        RECT 30.520 26.040 33.880 26.600 ;
        RECT 1.960 25.480 21.560 26.040 ;
        RECT 30.800 25.760 34.160 26.040 ;
        RECT 1.680 24.920 21.560 25.480 ;
        RECT 31.080 25.480 34.160 25.760 ;
        RECT 31.080 25.200 34.440 25.480 ;
        RECT 1.400 24.080 21.560 24.920 ;
        RECT 31.360 24.920 34.440 25.200 ;
        RECT 31.360 24.640 34.720 24.920 ;
        RECT 31.640 24.080 34.720 24.640 ;
        RECT 1.120 23.240 21.560 24.080 ;
        RECT 31.920 23.520 35.000 24.080 ;
        RECT 32.200 23.240 35.000 23.520 ;
        RECT 0.560 21.280 3.360 21.840 ;
        RECT 0.280 20.720 3.360 21.280 ;
        RECT 0.280 19.320 3.080 20.720 ;
        RECT 0.000 16.240 3.080 19.320 ;
        RECT 0.280 14.840 3.080 16.240 ;
        RECT 10.920 19.320 16.240 23.240 ;
        RECT 32.200 22.680 35.280 23.240 ;
        RECT 32.480 22.400 35.280 22.680 ;
        RECT 32.480 21.840 35.560 22.400 ;
        RECT 32.760 21.280 35.560 21.840 ;
        RECT 32.760 20.720 35.840 21.280 ;
        RECT 0.280 14.280 3.360 14.840 ;
        RECT 0.560 13.720 3.360 14.280 ;
        RECT 10.920 14.560 29.960 19.320 ;
        RECT 33.040 14.840 35.840 20.720 ;
        RECT 10.920 14.280 29.680 14.560 ;
        RECT 32.760 14.280 35.840 14.840 ;
        RECT 0.560 13.160 3.640 13.720 ;
        RECT 0.840 12.880 3.640 13.160 ;
        RECT 0.840 12.320 3.920 12.880 ;
        RECT 1.120 12.040 3.920 12.320 ;
        RECT 1.120 11.480 4.200 12.040 ;
        RECT 1.400 10.920 4.480 11.480 ;
        RECT 10.920 11.200 16.240 14.280 ;
        RECT 1.400 10.640 4.760 10.920 ;
        RECT 1.680 10.360 4.760 10.640 ;
        RECT 1.680 10.080 5.040 10.360 ;
        RECT 1.960 9.800 5.040 10.080 ;
        RECT 1.960 9.520 5.320 9.800 ;
        RECT 2.240 8.960 5.600 9.520 ;
        RECT 2.520 8.680 5.880 8.960 ;
        RECT 2.520 8.400 6.160 8.680 ;
        RECT 2.800 8.120 6.440 8.400 ;
        RECT 3.080 7.840 6.440 8.120 ;
        RECT 3.080 7.560 6.720 7.840 ;
        RECT 3.360 7.280 7.000 7.560 ;
        RECT 3.640 7.000 7.280 7.280 ;
        RECT 3.920 6.720 7.560 7.000 ;
        RECT 3.920 6.440 7.840 6.720 ;
        RECT 4.200 6.160 8.120 6.440 ;
        RECT 4.480 5.880 8.680 6.160 ;
        RECT 4.760 5.600 8.960 5.880 ;
        RECT 5.040 5.320 9.240 5.600 ;
        RECT 5.320 5.040 9.800 5.320 ;
        RECT 5.600 4.760 10.080 5.040 ;
        RECT 5.880 4.480 10.640 4.760 ;
        RECT 6.160 4.200 11.200 4.480 ;
        RECT 6.440 3.920 11.760 4.200 ;
        RECT 6.720 3.640 12.320 3.920 ;
        RECT 7.280 3.360 13.160 3.640 ;
        RECT 7.560 3.080 14.000 3.360 ;
        RECT 7.840 2.800 15.120 3.080 ;
        RECT 19.320 2.800 24.640 14.280 ;
        RECT 32.760 13.720 35.560 14.280 ;
        RECT 32.480 13.160 35.560 13.720 ;
        RECT 32.480 12.880 35.280 13.160 ;
        RECT 32.200 12.320 35.280 12.880 ;
        RECT 32.200 12.040 35.000 12.320 ;
        RECT 31.920 11.480 35.000 12.040 ;
        RECT 31.640 10.920 34.720 11.480 ;
        RECT 31.360 10.640 34.720 10.920 ;
        RECT 31.360 10.360 34.440 10.640 ;
        RECT 31.080 10.080 34.440 10.360 ;
        RECT 31.080 9.800 34.160 10.080 ;
        RECT 30.800 9.520 34.160 9.800 ;
        RECT 30.520 8.960 33.880 9.520 ;
        RECT 30.240 8.680 33.600 8.960 ;
        RECT 29.960 8.400 33.600 8.680 ;
        RECT 29.680 8.120 33.320 8.400 ;
        RECT 29.680 7.840 33.040 8.120 ;
        RECT 29.400 7.560 33.040 7.840 ;
        RECT 29.120 7.280 32.760 7.560 ;
        RECT 28.840 7.000 32.480 7.280 ;
        RECT 28.560 6.720 32.200 7.000 ;
        RECT 28.280 6.440 32.200 6.720 ;
        RECT 28.000 6.160 31.920 6.440 ;
        RECT 27.440 5.880 31.640 6.160 ;
        RECT 27.160 5.600 31.360 5.880 ;
        RECT 26.880 5.320 31.080 5.600 ;
        RECT 26.320 5.040 30.800 5.320 ;
        RECT 8.400 2.520 24.640 2.800 ;
        RECT 8.680 2.240 24.640 2.520 ;
        RECT 9.240 1.960 24.640 2.240 ;
        RECT 9.800 1.680 24.640 1.960 ;
        RECT 26.040 4.760 30.520 5.040 ;
        RECT 26.040 4.480 30.240 4.760 ;
        RECT 26.040 4.200 29.960 4.480 ;
        RECT 26.040 3.920 29.680 4.200 ;
        RECT 26.040 3.640 29.400 3.920 ;
        RECT 26.040 3.360 28.840 3.640 ;
        RECT 26.040 3.080 28.560 3.360 ;
        RECT 26.040 2.800 28.280 3.080 ;
        RECT 26.040 2.520 27.720 2.800 ;
        RECT 26.040 2.240 27.440 2.520 ;
        RECT 26.040 1.960 26.880 2.240 ;
        RECT 26.040 1.680 26.320 1.960 ;
        RECT 10.360 1.400 24.640 1.680 ;
        RECT 10.920 1.120 24.640 1.400 ;
        RECT 11.760 0.840 24.360 1.120 ;
        RECT 12.600 0.560 23.520 0.840 ;
        RECT 13.440 0.280 22.680 0.560 ;
        RECT 14.560 0.000 21.560 0.280 ;
  END
END ttlogo
END LIBRARY

